package ram_test_pkg;

	import uvm_pkg::*;
	
	`include "uvm_macros.svh"
	`include "seq_item.sv"
	`include "env_config.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "sequencer.sv"
	`include "src_agent.sv"
	`include "scoreboard.sv"

	`include "tb.sv"
	`include "base_seq.sv"
	
	`include "test.sv"
	 
endpackage
